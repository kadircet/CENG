`timescale 1ns / 1ps

module VBEncoder(input CLK,
			input [7:0] INT4,input [7:0] INT3, input [7:0] INT2, input [7:0] INT1,
            input START,
            output reg READY, 
			output reg [7:0] STREAM);

//Write your code below

endmodule